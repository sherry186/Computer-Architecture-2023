module ALU(data1_i, data2_i, ALUCtrl_i, data_o, Zero_o);
input signed [31:0] data1_i, data2_i;
input  [2:0]  ALUCtrl_i;
output [31:0] data_o;
output        Zero_o;

// TODO

endmodule
