module branch_predictor
(
    clk_i, 
    rst_i,

    update_i,
	result_i,
	predict_o
);
input clk_i, rst_i, update_i, result_i;
output predict_o;

// TODO

endmodule
